* C:\Users\HP\Desktop\208 project\Plant.sch

* Schematics Version 9.2
* Sun Aug 28 02:15:35 2022



** Analysis setup **
.tran 1u 500m 0 10u


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Plant.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
