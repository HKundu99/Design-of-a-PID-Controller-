* C:\Users\HP\Desktop\208 project\manual tuning.sch

* Schematics Version 9.2
* Sun Aug 28 09:25:12 2022



** Analysis setup **
.tran 100u 400m 0 100u


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "manual tuning.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
